** Profile: "SCHEMATIC1-phaseShift"  [ c:\users\amir\desktop\elec3\phaseshift\phaseshift-schematic1-phaseshift.sim ] 

** Creating circuit file "phaseshift-schematic1-phaseshift.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 10u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\phaseshift-SCHEMATIC1.net" 


.END
