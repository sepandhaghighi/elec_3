** Profile: "SCHEMATIC1-wien"  [ c:\users\amir\desktop\elec3\wien\wien-schematic1-wien.sim ] 

** Creating circuit file "wien-schematic1-wien.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 10u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\wien-SCHEMATIC1.net" 


.END
