** Profile: "SCHEMATIC1-noiseGenerator"  [ C:\USERS\AMIR\DESKTOP\ELEC3\noiseGenerator\noisegenerator-SCHEMATIC1-noiseGenerator.sim ] 

** Creating circuit file "noisegenerator-SCHEMATIC1-noiseGenerator.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\noisegenerator.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\noisegenerator-SCHEMATIC1.net" 


.END
